`define EQUATION0_ADDRESS_REG_OFFSET 8'h00
`define EQUATION1_ADDRESS_REG_OFFSET 8'h04
`define EQUATION2_ADDRESS_REG_OFFSET 8'h08
`define EQUATION3_ADDRESS_REG_OFFSET 8'h0C


`define CONTROL_REG_OFFSET          8'h10
`define CONTROL_REG_START_EQUATION0  0
`define CONTROL_REG_START_EQUATION1  1
`define CONTROL_REG_START_EQUATION2  2
`define CONTROL_REG_START_EQUATION3  3

`define CONTROL_REG_EQUATION_SELECT 3:0
`define CONTROL_REG_STOP_EQUATION   4
`define CONTROL_REG_BEGIN_EQUATION  5
`define CONTROL_REG_SIGNED_DATA     6
`define CONTROL_EQUATION_EQUATION   31:24

`define STATUS_REG_OFFSET           8'h14
`define STATUS_REG_ACTIVE           0

//
// Equation Structure
//
`define EQUATION_CONTROL_OFFSET       8'h00
`define EQUATION_STATUS_OFFSET        8'h04
`define EQUATION_NEXT_ADDRESS_OFFSET  8'h08
`define EQUATION_RESERVED0_OFFSET     8'h0C
`define EQUATION_X_VECTOR_OFFSET      8'h10
`define EQUATION_Y_VECTOR_OFFSET      8'h30
`define EQUATION_Z_VECTOR_OFFSET      8'h50
`define EQUATION_RESULT_VECTOR_OFFSET 8'h70

`define EQUATION_CONTROL_SELECT_NONE  8'h00
`define EQUATION_CONTROL_SELECT_SUM   8'h01
