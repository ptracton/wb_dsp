`define DAQ_CONTROL_REG_OFFSET      8'h0

`define DAQ_CHANNEL0_ADDRESS_OFFSET 8'h10
`define DAQ_CHANNEL1_ADDRESS_OFFSET 8'h20
`define DAQ_CHANNEL2_ADDRESS_OFFSET 8'h40
`define DAQ_CHANNEL3_ADDRESS_OFFSET 8'h80

/**
 Vector Structure
 **/
`define VECTOR_CONTROL_OFFSET        8'h00
`define VECTOR_STATUS_OFFSET         8'h04
`define VECTOR_START_ADDRESS_OFFSET  8'h08
`define VECTOR_END_ADDRESS_OFFSET    8'h0C 
`define VECTOR_READ_POINTER_OFFSET   8'h10
`define VECTOR_WRITE_POINTER_OFFSET  8'h14
`define VECTOR_RESERVED0_OFFSET      8'h18
`define VECTOR_RESERVED1_OFFSET      8'h1C


