`define DAQ_CONTROL_REG_OFFSET      8'h0

`define DAQ_CHANNEL0_ADDRESS_OFFSET 8'h10
`define DAQ_CHANNEL0_CONTROL_OFFSET 8'h14
`define DAQ_CHANNEL0_STATUS_OFFSET  8'h18

`define DAQ_CHANNEL1_ADDRESS_OFFSET 8'h20
`define DAQ_CHANNEL1_CONTROL_OFFSET 8'h24
`define DAQ_CHANNEL1_STATUS_OFFSET  8'h28

`define DAQ_CHANNEL2_ADDRESS_OFFSET 8'h30
`define DAQ_CHANNEL2_CONTROL_OFFSET 8'h34
`define DAQ_CHANNEL2_STATUS_OFFSET  8'h38

`define DAQ_CHANNEL3_ADDRESS_OFFSET 8'h40
`define DAQ_CHANNEL3_CONTROL_OFFSET 8'h44
`define DAQ_CHANNEL3_STATUS_OFFSET  8'h48

/**
 DAQ Channel Control Register Bits
 **/
`define DAQ_CHANNEL_ENABLE_OFFSET         0
`define DAQ_CHANNEL_SIGNED_OFFSET         1
`define DAQ_CHANNEL_ADC_CLK_SPEED_OFFSET  2  // 3 bits wide
`define DAQ_CHANNEL_ADC_DATA_WIDTH_OFFSET 5  // 3 bits wide
`define DAQ_CHANNEL_DECIMATOR_SELECT      8  // 2 bits wide
`define DAQ_CHANNEL_FIFO_SAMPLES          10 // 6 bits wide
`define DAQ_CHANNEL_SAMPLES_PER_EQUATION  16 // 8 bits wide

`define DAQ_CHANNEL_ENABLE 1 << `DAQ_CHANNEL_ENABLE_OFFSET
`define DAQ_CHANNEL_SIGNED 1 << `DAQ_CHANNEL_SIGNED_OFFSET


/**
 Vector Structure
 **/
`define VECTOR_CONTROL_OFFSET        8'h00
`define VECTOR_STATUS_OFFSET         8'h04
`define VECTOR_START_ADDRESS_OFFSET  8'h08
`define VECTOR_END_ADDRESS_OFFSET    8'h0C 
`define VECTOR_READ_POINTER_OFFSET   8'h10
`define VECTOR_WRITE_POINTER_OFFSET  8'h14
`define VECTOR_RESERVED0_OFFSET      8'h18
`define VECTOR_RESERVED1_OFFSET      8'h1C


