`define EQUATION_ADDRESS_REG_OFFSET 4'h0


`define CONTROL_REG_OFFSET          4'h4
`define CONTROL_REG_START_EQUATION  0
`define CONTROL_REG_STOP_EQUATION   1
`define CONTROL_EQUATION_EQUATION   31:24

`define STATUS_REG_OFFSET           4'h8
`define STATUS_REG_ACTIVE           0
